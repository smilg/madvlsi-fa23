magic
tech sky130A
timestamp 1695745633
<< nwell >>
rect 45 5 385 505
<< nmos >>
rect 115 -525 130 -140
rect 170 -240 185 -140
rect 235 -240 250 -140
rect 300 -240 315 -140
rect 170 -525 185 -425
rect 235 -525 250 -425
rect 300 -525 315 -425
<< pmos >>
rect 115 310 130 410
rect 180 310 195 410
rect 115 25 130 125
rect 180 25 195 125
rect 245 25 260 410
rect 300 310 315 410
rect 300 25 315 125
<< ndiff >>
rect 65 -155 115 -140
rect 65 -510 80 -155
rect 100 -510 115 -155
rect 65 -525 115 -510
rect 130 -240 170 -140
rect 185 -155 235 -140
rect 185 -225 200 -155
rect 220 -225 235 -155
rect 185 -240 235 -225
rect 250 -155 300 -140
rect 250 -225 265 -155
rect 285 -225 300 -155
rect 250 -240 300 -225
rect 315 -155 365 -140
rect 315 -225 330 -155
rect 350 -225 365 -155
rect 315 -240 365 -225
rect 130 -425 155 -240
rect 130 -525 170 -425
rect 185 -440 235 -425
rect 185 -510 200 -440
rect 220 -510 235 -440
rect 185 -525 235 -510
rect 250 -440 300 -425
rect 250 -510 265 -440
rect 285 -510 300 -440
rect 250 -525 300 -510
rect 315 -440 365 -425
rect 315 -510 330 -440
rect 350 -510 365 -440
rect 315 -525 365 -510
<< pdiff >>
rect 65 395 115 410
rect 65 325 80 395
rect 100 325 115 395
rect 65 310 115 325
rect 130 395 180 410
rect 130 325 145 395
rect 165 325 180 395
rect 130 310 180 325
rect 195 395 245 410
rect 195 325 210 395
rect 230 325 245 395
rect 195 310 245 325
rect 220 125 245 310
rect 65 110 115 125
rect 65 40 80 110
rect 100 40 115 110
rect 65 25 115 40
rect 130 110 180 125
rect 130 40 145 110
rect 165 40 180 110
rect 130 25 180 40
rect 195 110 245 125
rect 195 40 210 110
rect 230 40 245 110
rect 195 25 245 40
rect 260 310 300 410
rect 315 395 365 410
rect 315 325 330 395
rect 350 325 365 395
rect 315 310 365 325
rect 260 125 285 310
rect 260 25 300 125
rect 315 110 365 125
rect 315 40 330 110
rect 350 40 365 110
rect 315 25 365 40
<< ndiffc >>
rect 80 -510 100 -155
rect 200 -225 220 -155
rect 265 -225 285 -155
rect 330 -225 350 -155
rect 200 -510 220 -440
rect 265 -510 285 -440
rect 330 -510 350 -440
<< pdiffc >>
rect 80 325 100 395
rect 145 325 165 395
rect 210 325 230 395
rect 80 40 100 110
rect 145 40 165 110
rect 210 40 230 110
rect 330 325 350 395
rect 330 40 350 110
<< psubdiff >>
rect 265 -570 365 -555
rect 265 -590 280 -570
rect 350 -590 365 -570
rect 265 -605 365 -590
<< nsubdiff >>
rect 170 472 270 487
rect 170 452 185 472
rect 255 452 270 472
rect 170 437 270 452
<< psubdiffcont >>
rect 280 -590 350 -570
<< nsubdiffcont >>
rect 185 452 255 472
<< poly >>
rect 115 410 130 425
rect 180 410 195 425
rect 245 410 260 425
rect 300 410 315 425
rect 115 295 130 310
rect 70 280 130 295
rect 70 155 85 280
rect 180 255 195 310
rect 106 245 195 255
rect 106 225 116 245
rect 136 240 195 245
rect 136 225 146 240
rect 106 215 146 225
rect 165 190 205 200
rect 165 170 175 190
rect 195 170 205 190
rect 165 160 205 170
rect 70 140 130 155
rect 115 125 130 140
rect 180 125 195 160
rect 300 295 315 310
rect 300 285 365 295
rect 300 280 335 285
rect 325 265 335 280
rect 355 265 365 285
rect 325 255 365 265
rect 300 125 315 140
rect 115 -140 130 25
rect 180 -35 195 25
rect 245 10 260 25
rect 235 -5 260 10
rect 170 -45 210 -35
rect 170 -65 180 -45
rect 200 -65 210 -45
rect 170 -75 210 -65
rect 170 -140 185 -125
rect 235 -140 250 -5
rect 300 -20 315 25
rect 275 -30 315 -20
rect 275 -50 285 -30
rect 305 -50 315 -30
rect 275 -60 315 -50
rect 315 -95 355 -85
rect 315 -105 325 -95
rect 300 -115 325 -105
rect 345 -115 355 -95
rect 300 -125 355 -115
rect 300 -140 315 -125
rect 170 -295 185 -240
rect 235 -255 250 -240
rect 300 -255 315 -240
rect 235 -270 255 -255
rect 300 -265 360 -255
rect 300 -270 330 -265
rect 170 -305 210 -295
rect 170 -325 180 -305
rect 200 -325 210 -305
rect 170 -335 210 -325
rect 173 -367 213 -357
rect 173 -387 183 -367
rect 203 -387 213 -367
rect 173 -397 213 -387
rect 240 -395 255 -270
rect 320 -285 330 -270
rect 350 -285 360 -265
rect 320 -295 360 -285
rect 280 -330 320 -320
rect 280 -350 290 -330
rect 310 -350 320 -330
rect 280 -360 320 -350
rect 170 -410 190 -397
rect 235 -410 255 -395
rect 170 -425 185 -410
rect 235 -425 250 -410
rect 300 -425 315 -360
rect 115 -630 130 -525
rect 170 -540 185 -525
rect 235 -630 250 -525
rect 300 -540 315 -525
rect 90 -640 130 -630
rect 90 -660 100 -640
rect 120 -660 130 -640
rect 90 -670 130 -660
rect 210 -640 250 -630
rect 210 -660 220 -640
rect 240 -660 250 -640
rect 210 -670 250 -660
<< polycont >>
rect 116 225 136 245
rect 175 170 195 190
rect 335 265 355 285
rect 180 -65 200 -45
rect 285 -50 305 -30
rect 325 -115 345 -95
rect 180 -325 200 -305
rect 183 -387 203 -367
rect 330 -285 350 -265
rect 290 -350 310 -330
rect 100 -660 120 -640
rect 220 -660 240 -640
<< locali >>
rect 175 472 265 482
rect 175 452 185 472
rect 255 452 265 472
rect 175 442 265 452
rect 70 395 110 405
rect 70 335 80 395
rect 45 325 80 335
rect 100 325 110 395
rect 45 315 110 325
rect 135 395 175 405
rect 135 325 145 395
rect 165 325 175 395
rect 135 315 175 325
rect 200 395 240 442
rect 200 325 210 395
rect 230 325 240 395
rect 320 395 360 405
rect 320 335 330 395
rect 200 315 240 325
rect 265 325 330 335
rect 350 335 360 395
rect 350 325 385 335
rect 265 315 385 325
rect 155 295 175 315
rect 155 275 195 295
rect 106 245 146 255
rect 106 225 116 245
rect 136 225 146 245
rect 106 215 146 225
rect 115 160 135 215
rect 175 200 195 275
rect 165 190 205 200
rect 165 170 175 190
rect 195 170 205 190
rect 165 160 205 170
rect 115 140 145 160
rect 128 120 155 140
rect 45 110 110 120
rect 45 100 80 110
rect 70 40 80 100
rect 100 40 110 110
rect 70 30 110 40
rect 135 110 175 120
rect 135 40 145 110
rect 165 40 175 110
rect 135 30 175 40
rect 200 110 240 120
rect 200 40 210 110
rect 230 40 240 110
rect 200 30 240 40
rect 135 5 155 30
rect 115 -15 155 5
rect 115 -100 135 -15
rect 265 -20 285 315
rect 325 285 365 295
rect 325 265 335 285
rect 355 265 365 285
rect 325 255 365 265
rect 325 120 345 255
rect 320 110 385 120
rect 320 40 330 110
rect 350 100 385 110
rect 350 40 360 100
rect 320 30 360 40
rect 265 -30 315 -20
rect 265 -35 285 -30
rect 170 -45 210 -35
rect 170 -65 180 -45
rect 200 -65 210 -45
rect 170 -75 210 -65
rect 115 -120 155 -100
rect 70 -155 110 -145
rect 70 -510 80 -155
rect 100 -510 110 -155
rect 135 -295 155 -120
rect 190 -145 210 -75
rect 275 -50 285 -35
rect 305 -50 315 -30
rect 275 -60 315 -50
rect 275 -145 295 -60
rect 335 -85 355 30
rect 315 -95 355 -85
rect 315 -115 325 -95
rect 345 -115 355 -95
rect 315 -125 355 -115
rect 190 -155 230 -145
rect 190 -225 200 -155
rect 220 -225 230 -155
rect 190 -235 230 -225
rect 255 -155 295 -145
rect 255 -225 265 -155
rect 285 -225 295 -155
rect 255 -235 295 -225
rect 320 -155 360 -145
rect 320 -225 330 -155
rect 350 -225 360 -155
rect 320 -235 360 -225
rect 210 -255 230 -235
rect 210 -275 250 -255
rect 135 -305 210 -295
rect 135 -325 180 -305
rect 200 -325 210 -305
rect 135 -335 210 -325
rect 135 -430 155 -335
rect 230 -355 250 -275
rect 275 -320 295 -235
rect 320 -265 360 -255
rect 320 -285 330 -265
rect 350 -285 360 -265
rect 320 -295 360 -285
rect 275 -330 320 -320
rect 210 -357 250 -355
rect 173 -367 250 -357
rect 280 -350 290 -330
rect 310 -350 320 -330
rect 280 -360 320 -350
rect 173 -387 183 -367
rect 203 -375 250 -367
rect 203 -387 213 -375
rect 173 -397 213 -387
rect 340 -390 360 -295
rect 275 -410 360 -390
rect 275 -430 295 -410
rect 135 -440 230 -430
rect 135 -450 200 -440
rect 70 -520 110 -510
rect 190 -510 200 -450
rect 220 -510 230 -440
rect 190 -520 230 -510
rect 255 -440 295 -430
rect 255 -510 265 -440
rect 285 -510 295 -440
rect 255 -520 295 -510
rect 320 -440 360 -430
rect 320 -510 330 -440
rect 350 -510 360 -440
rect 320 -560 360 -510
rect 270 -570 360 -560
rect 270 -590 280 -570
rect 350 -590 360 -570
rect 270 -600 360 -590
rect 90 -640 130 -630
rect 90 -660 100 -640
rect 120 -660 130 -640
rect 90 -670 130 -660
rect 210 -640 250 -630
rect 210 -660 220 -640
rect 240 -660 250 -640
rect 210 -670 250 -660
<< viali >>
rect 185 452 255 472
rect 210 325 230 395
rect 210 40 230 110
rect 80 -510 100 -155
rect 330 -225 350 -155
rect 330 -510 350 -440
rect 280 -590 350 -570
rect 100 -660 120 -640
rect 220 -660 240 -640
<< metal1 >>
rect 45 472 385 490
rect 45 452 185 472
rect 255 452 385 472
rect 45 395 385 452
rect 45 325 210 395
rect 230 325 385 395
rect 45 110 385 325
rect 45 40 210 110
rect 230 40 385 110
rect 45 25 385 40
rect 280 -25 300 25
rect 45 -155 385 -140
rect 45 -510 80 -155
rect 100 -225 330 -155
rect 350 -225 385 -155
rect 100 -440 385 -225
rect 100 -510 330 -440
rect 350 -510 385 -440
rect 45 -570 385 -510
rect 45 -590 280 -570
rect 350 -590 385 -570
rect 45 -600 385 -590
rect 45 -640 385 -630
rect 45 -660 100 -640
rect 120 -660 220 -640
rect 240 -660 385 -640
rect 45 -670 385 -660
<< labels >>
rlabel metal1 45 465 45 465 7 VP
port 6 w
rlabel locali 45 325 45 325 7 D
port 1 w
rlabel locali 45 110 45 110 7 Db
port 2 w
rlabel metal1 45 -580 45 -580 7 VN
port 7 w
rlabel metal1 45 -650 45 -650 7 CLK
port 3 w
rlabel locali 385 325 385 325 3 Q
port 4 e
rlabel locali 385 110 385 110 3 Qb
port 5 e
<< end >>
