magic
tech sky130A
timestamp 1694461190
<< nwell >>
rect -120 135 150 275
<< nmos >>
rect 0 0 15 100
rect 65 0 80 100
<< pmos >>
rect 0 155 15 255
rect 65 155 80 255
<< ndiff >>
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 0 65 100
rect 80 85 130 100
rect 80 15 95 85
rect 115 15 130 85
rect 80 0 130 15
<< pdiff >>
rect -50 240 0 255
rect -50 170 -35 240
rect -15 170 0 240
rect -50 155 0 170
rect 15 240 65 255
rect 15 170 30 240
rect 50 170 65 240
rect 15 155 65 170
rect 80 240 130 255
rect 80 170 95 240
rect 115 170 130 240
rect 80 155 130 170
<< ndiffc >>
rect -35 15 -15 85
rect 95 15 115 85
<< pdiffc >>
rect -35 170 -15 240
rect 30 170 50 240
rect 95 170 115 240
<< psubdiff >>
rect -100 85 -50 100
rect -100 15 -85 85
rect -65 15 -50 85
rect -100 0 -50 15
<< nsubdiff >>
rect -100 240 -50 255
rect -100 170 -85 240
rect -65 170 -50 240
rect -100 155 -50 170
<< psubdiffcont >>
rect -85 15 -65 85
<< nsubdiffcont >>
rect -85 170 -65 240
<< poly >>
rect 0 255 15 270
rect 65 255 80 270
rect 0 100 15 155
rect 65 100 80 155
rect 0 -15 15 0
rect 65 -15 80 0
rect -25 -25 15 -15
rect -25 -45 -15 -25
rect 5 -45 15 -25
rect -25 -55 15 -45
rect 40 -25 80 -15
rect 40 -45 50 -25
rect 70 -45 80 -25
rect 40 -55 80 -45
<< polycont >>
rect -15 -45 5 -25
rect 50 -45 70 -25
<< locali >>
rect -95 240 -5 250
rect -95 170 -85 240
rect -65 170 -35 240
rect -15 170 -5 240
rect -95 160 -5 170
rect 20 240 60 250
rect 20 170 30 240
rect 50 170 60 240
rect 20 160 60 170
rect 85 240 125 250
rect 85 170 95 240
rect 115 170 125 240
rect 85 160 125 170
rect 40 140 60 160
rect 40 120 105 140
rect 85 95 105 120
rect -95 85 -5 95
rect -95 15 -85 85
rect -65 15 -35 85
rect -15 15 -5 85
rect -95 5 -5 15
rect 85 85 125 95
rect 85 15 95 85
rect 115 15 125 85
rect 85 5 125 15
rect 105 -15 125 5
rect -120 -25 15 -15
rect -120 -35 -15 -25
rect -25 -45 -15 -35
rect 5 -45 15 -25
rect -25 -55 15 -45
rect 40 -25 80 -15
rect 40 -45 50 -25
rect 70 -45 80 -25
rect 105 -35 150 -15
rect 40 -55 80 -45
rect -120 -75 -45 -55
rect 40 -75 60 -55
rect -65 -95 60 -75
<< viali >>
rect -85 170 -65 240
rect -35 170 -15 240
rect 95 170 115 240
rect -85 15 -65 85
rect -35 15 -15 85
<< metal1 >>
rect -120 240 150 250
rect -120 170 -85 240
rect -65 170 -35 240
rect -15 170 95 240
rect 115 170 150 240
rect -120 160 150 170
rect -120 85 150 95
rect -120 15 -85 85
rect -65 15 -35 85
rect -15 15 150 85
rect -120 5 150 15
<< labels >>
rlabel locali -120 -25 -120 -25 7 A
port 1 w
rlabel locali -120 -65 -120 -65 7 B
port 2 w
rlabel locali 150 -25 150 -25 3 Y
port 3 e
rlabel metal1 -120 205 -120 205 7 VP
port 4 w
rlabel metal1 -120 50 -120 50 7 VN
port 5 w
<< end >>
