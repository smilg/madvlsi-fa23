magic
tech sky130A
timestamp 1694461552
<< locali >>
rect 0 60 25 80
rect 450 60 475 80
rect 0 20 25 40
<< metal1 >>
rect 0 255 25 345
rect 0 100 25 190
use inverter  inverter_0
timestamp 1694458850
transform 1 0 390 0 1 95
box -120 -55 85 275
use NAND2  NAND2_0
timestamp 1694461190
transform 1 0 120 0 1 95
box -120 -95 150 275
<< labels >>
rlabel locali 0 70 0 70 7 A
rlabel locali 0 30 0 30 7 B
rlabel metal1 0 300 0 300 7 VP
rlabel metal1 0 145 0 145 7 VN
rlabel locali 475 70 475 70 3 Y
<< end >>
